----------------------------------
-- Engineer: Eros Garcia Arroyo --
----------------------------------

---------------
-- Libraries --
---------------
library ieee;
use ieee.std_logic_1164.all;

-------------
-- Package --
-------------
package pkg_digital_effects is

  component efecto_es is
    generic(
      g_width : integer := 12 --Ancho del bus
    ); 
    port( 
      clk        : in std_logic;
      reset_n    : in std_logic; 
      enable_in  : in std_logic;
      l_data_in  : in std_logic_vector(g_width-1 downto 0);                        
      r_data_in  : in std_logic_vector(g_width-1 downto 0);                          
      l_data_out : out std_logic_vector(g_width-1 downto 0);                           
      r_data_out : out std_logic_vector(g_width-1 downto 0) 
    );
  end component;

  component efecto_delay is
    generic(
      n       : integer := 4000;
      g_width : integer := 12);
    port( 
      clk        : in std_logic;   
      reset_n    : in std_logic;   
      enable_in  : in std_logic;   
      l_data_in  : in std_logic_vector(g_width-1 downto 0);             
      r_data_in  : in std_logic_vector(g_width-1 downto 0);                             
      l_data_out : out std_logic_vector(g_width-1 downto 0);                        
      r_data_out : out std_logic_vector(g_width-1 downto 0)
    ); 
  end component;

  component efecto_chorus is
    generic(
      n       : integer := 1000;
      g_width : integer := 12);
    port( 
      clk        : in std_logic;   
      reset_n    : in std_logic;   
      enable_in  : in std_logic;   
      l_data_in  : in std_logic_vector(g_width-1 downto 0);             
      r_data_in  : in std_logic_vector(g_width-1 downto 0);                             
      l_data_out : out std_logic_vector(g_width-1 downto 0);                        
      r_data_out : out std_logic_vector(g_width-1 downto 0)
    ); 
  end component;

  component efecto_vibrato is
    generic(
      n       : integer := 500;
      g_width : integer := 12 
    );
    port( 
      clk        : in std_logic;                                         
      reset_n    : in std_logic;
      enable_in  : in std_logic; 
      l_data_in  : in std_logic_vector(g_width-1 downto 0);                         
      r_data_in  : in std_logic_vector(g_width-1 downto 0);                           
      l_data_out : out std_logic_vector(g_width-1 downto 0);                            
      r_data_out : out std_logic_vector(g_width-1 downto 0) 
  ); 
  end component;

  component efecto_reverb is
    generic(
      n       : integer := 500;
      g_width : integer := 12 
    );
    port( 
      clk        : in std_logic; 
      reset_n    : in std_logic; 
      enable_in  : in std_logic; 
      l_data_in  : in std_logic_vector(g_width-1 downto 0);                      
      r_data_in  : in std_logic_vector(g_width-1 downto 0);                        
      l_data_out : out std_logic_vector(g_width-1 downto 0);                         
      r_data_out : out std_logic_vector(g_width-1 downto 0) 
    ); 
  end component;

  component efecto_eco is
    generic(
      n       : integer := 5000;
      g_width : integer := 12 
    );
    port( 
      clk        : in std_logic; 
      reset_n    : in std_logic; 
      enable_in  : in std_logic; 
      l_data_in  : in std_logic_vector(g_width-1 downto 0);                      
      r_data_in  : in std_logic_vector(g_width-1 downto 0);                        
      l_data_out : out std_logic_vector(g_width-1 downto 0);                         
      r_data_out : out std_logic_vector(g_width-1 downto 0) 
    ); 
  end component;

  component efecto_compressor is
    generic(
      g_width : integer := 12 
      );
    port ( 
      clk        : in std_logic;   
      reset_n    : in std_logic;   
      enable_in  : in std_logic;   
      l_data_in  : in std_logic_vector(g_width-1 downto 0);             
      r_data_in  : in std_logic_vector(g_width-1 downto 0);                             
      l_data_out : out std_logic_vector(g_width-1 downto 0);                        
      r_data_out : out std_logic_vector(g_width-1 downto 0)
  );
  end component;

  component efecto_overdrive is
    generic(
      g_width : integer := 12 
      );
    port ( 
      clk        : in std_logic;    
      reset_n    : in std_logic;    
      enable_in  : in std_logic;    
      l_data_in  : in std_logic_vector(g_width-1 downto 0);             
      r_data_in  : in std_logic_vector(g_width-1 downto 0);                             
      l_data_out : out std_logic_vector(g_width-1 downto 0);                        
      r_data_out : out std_logic_vector(g_width-1 downto 0)
    );
  end component;

component EfectoLOOPER is
GENERIC(
    d_width         : INTEGER := 12;
    d_deep          : INTEGER := 19
    );
Port ( 
    clk                   : in STD_LOGIC;
    reset_n               : in STD_LOGIC;
    SW13                  : in STD_LOGIC;
    enable_in             : IN STD_LOGIC;
    SW5                   : IN STD_LOGIC;
    SW6                   : IN STD_LOGIC;
    l_data_in             : in STD_LOGIC_VECTOR (d_width-1  downto 0); -- STD_LOGIC;
    l_data_out            : out STD_LOGIC_VECTOR (d_width-1  downto 0);
    r_data_in             : in STD_LOGIC_VECTOR (d_width-1  downto 0); -- STD_LOGIC;
    r_data_out            : out STD_LOGIC_VECTOR (d_width-1  downto 0);
    enable_out            : out STD_LOGIC
);
end component;

component EfectoBANKFILTER is
GENERIC(
    d_width         :  INTEGER := 12);
Port ( 
    clk                   : in STD_LOGIC;
    reset_n               : in STD_LOGIC;
    enable_in             : in STD_LOGIC;
    SW14                  : IN STD_LOGIC; --Switch de control para el tipo de filtro
    l_data_in             : in STD_LOGIC_VECTOR (d_width-1  downto 0); -- STD_LOGIC;
    l_data_out            : out STD_LOGIC_VECTOR (d_width-1  downto 0);
    r_data_in             : in STD_LOGIC_VECTOR (d_width-1  downto 0); -- STD_LOGIC;
    r_data_out            : out STD_LOGIC_VECTOR (d_width-1  downto 0);
    enable_out            : out STD_LOGIC  
); 
end component;

  component efecto_config_reverb is
    generic(
      n1      : integer := 1500;
      g_width : integer := 12); 
    port( 
      clk        : in std_logic;
      reset_n    : in std_logic;
      enable_in  : in std_logic;
      BTNC       : in std_logic;
      BTNL       : in std_logic;
      BTND       : in std_logic;
      BTNR       : in std_logic;
      l_data_in  : in std_logic_vector(g_width-1 downto 0);                         
      r_data_in  : in std_logic_vector(g_width-1 downto 0);                           
      l_data_out : out std_logic_vector(g_width-1 downto 0);                            
      r_data_out : out std_logic_vector(g_width-1 downto 0) 
    ); 
  end component;

    
end pkg_digital_effects;